module counter (
input a,b
output q
);


endmodule