module counter (
input a,b
output q
// hola esto es un comentario 
);
reg temp;
asign q = temp;  
always @ a begin
    temp=temp+1:
end

endmodule